module adder_AXI_tb ();

    timeunit 1ns/1ps;

    localparam WIDTH  = 8;
    
endmodule